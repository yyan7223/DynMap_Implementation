
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_runOne.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_runOne.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_runOne.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_runOne.grp_Reset_fu_334.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_runOne.grp_Reset_fu_334.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_692_8_VITIS_LOOP_693_9_fu_197.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_692_8_VITIS_LOOP_693_9_fu_197.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_692_8_VITIS_LOOP_693_9_fu_197.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_704_13_fu_209.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_704_13_fu_209.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_704_13_fu_209.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_707_14_fu_215.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_707_14_fu_215.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_707_14_fu_215.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_710_15_fu_221.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_710_15_fu_221.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_710_15_fu_221.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_713_16_fu_227.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_713_16_fu_227.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_713_16_fu_227.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_716_17_fu_233.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_716_17_fu_233.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_716_17_fu_233.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_624_6_fu_430.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_624_6_fu_430.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_624_6_fu_430.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_453_4_fu_530.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_453_4_fu_530.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_453_4_fu_530.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_ready;
    assign module_intf_23.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_done;
    assign module_intf_23.ap_continue = 1'b1;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_577_16_fu_575.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_577_16_fu_575.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_577_16_fu_575.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_518_12_fu_584.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_518_12_fu_584.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_518_12_fu_584.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_480_7_fu_592.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_480_7_fu_592.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_480_7_fu_592.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_388_2_fu_482.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_388_2_fu_482.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_388_2_fu_482.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_ready;
    assign module_intf_30.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_done;
    assign module_intf_30.ap_continue = 1'b1;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ready;
    assign module_intf_31.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_done;
    assign module_intf_31.ap_continue = 1'b1;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ready;
    assign module_intf_37.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_done;
    assign module_intf_37.ap_continue = 1'b1;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_249_4_fu_402.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_249_4_fu_402.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_249_4_fu_402.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ready;
    assign module_intf_41.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_done;
    assign module_intf_41.ap_continue = 1'b1;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ready;
    assign module_intf_49.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_done;
    assign module_intf_49.ap_continue = 1'b1;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_start;
    assign module_intf_50.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ready;
    assign module_intf_50.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_done;
    assign module_intf_50.ap_continue = 1'b1;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;

    pp_loop_intf #(15) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_state1;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_state15;
    assign pp_loop_intf_1.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_1.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_state16;
    assign pp_loop_intf_1.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_enable_reg_pp0_iter1;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.quit_at_end = 1'b1;
    assign pp_loop_intf_1.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_354_4_fu_700.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(15) pp_loop_monitor_1;
    seq_loop_intf#(59) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_runOne.ap_ST_fsm_state54;
    assign seq_loop_intf_1.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.pre_loop_state1 = 59'h0;
    assign seq_loop_intf_1.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.pre_loop_state2 = 59'h0;
    assign seq_loop_intf_1.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_runOne.ap_ST_fsm_state1;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 59'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state2 = 59'h0;
    assign seq_loop_intf_1.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.post_loop_state3 = 59'h0;
    assign seq_loop_intf_1.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_runOne.ap_ST_fsm_state55;
    assign seq_loop_intf_1.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.quit_loop_state1 = 59'h0;
    assign seq_loop_intf_1.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state2 = 59'h0;
    assign seq_loop_intf_1.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.cur_state = AESL_inst_runOne.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_runOne.ap_ST_fsm_state55;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_runOne.ap_ST_fsm_state59;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(59) seq_loop_monitor_1;
    seq_loop_intf#(7) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state2;
    assign seq_loop_intf_2.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_2.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.pre_loop_state2 = 7'h0;
    assign seq_loop_intf_2.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state4;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 7'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.post_loop_state2 = 7'h0;
    assign seq_loop_intf_2.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.post_loop_state3 = 7'h0;
    assign seq_loop_intf_2.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state3;
    assign seq_loop_intf_2.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_2.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state2 = 7'h0;
    assign seq_loop_intf_2.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.cur_state = AESL_inst_runOne.grp_Reset_fu_334.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state3;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state3;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b1;
    assign seq_loop_intf_2.one_state_block = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state3_blk;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(7) seq_loop_monitor_2;
    seq_loop_intf#(7) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state3;
    assign seq_loop_intf_3.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_3.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.pre_loop_state2 = 7'h0;
    assign seq_loop_intf_3.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state5;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 7'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state2 = 7'h0;
    assign seq_loop_intf_3.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.post_loop_state3 = 7'h0;
    assign seq_loop_intf_3.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state4;
    assign seq_loop_intf_3.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_3.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state2 = 7'h0;
    assign seq_loop_intf_3.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.cur_state = AESL_inst_runOne.grp_Reset_fu_334.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state4;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state4;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b1;
    assign seq_loop_intf_3.one_state_block = AESL_inst_runOne.grp_Reset_fu_334.ap_ST_fsm_state4_blk;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(7) seq_loop_monitor_3;
    seq_loop_intf#(30) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state5;
    assign seq_loop_intf_4.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.pre_loop_state1 = 30'h0;
    assign seq_loop_intf_4.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.pre_loop_state2 = 30'h0;
    assign seq_loop_intf_4.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state16;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state18;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_4.post_loop_state2 = 30'h0;
    assign seq_loop_intf_4.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.post_loop_state3 = 30'h0;
    assign seq_loop_intf_4.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state6;
    assign seq_loop_intf_4.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.quit_loop_state1 = 30'h0;
    assign seq_loop_intf_4.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state2 = 30'h0;
    assign seq_loop_intf_4.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state6;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state14;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(30) seq_loop_monitor_4;
    seq_loop_intf#(30) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state17;
    assign seq_loop_intf_5.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.pre_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state25;
    assign seq_loop_intf_5.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_5.pre_loop_state2 = 30'h0;
    assign seq_loop_intf_5.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state29;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = 30'h0;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.post_loop_state2 = 30'h0;
    assign seq_loop_intf_5.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_5.post_loop_state3 = 30'h0;
    assign seq_loop_intf_5.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state26;
    assign seq_loop_intf_5.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.quit_loop_state1 = 30'h0;
    assign seq_loop_intf_5.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state2 = 30'h0;
    assign seq_loop_intf_5.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_5.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state26;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state28;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(30) seq_loop_monitor_5;
    seq_loop_intf#(30) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state1;
    assign seq_loop_intf_6.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.pre_loop_state1 = 30'h0;
    assign seq_loop_intf_6.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.pre_loop_state2 = 30'h0;
    assign seq_loop_intf_6.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state30;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 30'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.post_loop_state2 = 30'h0;
    assign seq_loop_intf_6.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_6.post_loop_state3 = 30'h0;
    assign seq_loop_intf_6.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state3;
    assign seq_loop_intf_6.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.quit_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state29;
    assign seq_loop_intf_6.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_6.quit_loop_state2 = 30'h0;
    assign seq_loop_intf_6.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_6.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state2;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.ap_ST_fsm_state29;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(30) seq_loop_monitor_6;
    seq_loop_intf#(5) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state1;
    assign seq_loop_intf_7.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_7.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_7.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state4;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state5;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_7.post_loop_state2 = 5'h0;
    assign seq_loop_intf_7.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_7.post_loop_state3 = 5'h0;
    assign seq_loop_intf_7.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state3;
    assign seq_loop_intf_7.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_7.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_7.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_7.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state2;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_601_2_fu_403.ap_ST_fsm_state3;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(5) seq_loop_monitor_7;
    seq_loop_intf#(5) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state1;
    assign seq_loop_intf_8.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_8.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_8.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state4;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state5;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_8.post_loop_state2 = 5'h0;
    assign seq_loop_intf_8.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_8.post_loop_state3 = 5'h0;
    assign seq_loop_intf_8.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state3;
    assign seq_loop_intf_8.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_8.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_8.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_8.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_611_4_fu_411.ap_ST_fsm_state3;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(5) seq_loop_monitor_8;
    seq_loop_intf#(5) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state1;
    assign seq_loop_intf_9.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_9.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_9.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state4;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state5;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_9.post_loop_state2 = 5'h0;
    assign seq_loop_intf_9.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_9.post_loop_state3 = 5'h0;
    assign seq_loop_intf_9.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state3;
    assign seq_loop_intf_9.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_9.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_9.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_9.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state2;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_618_5_fu_422.ap_ST_fsm_state3;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(5) seq_loop_monitor_9;
    seq_loop_intf#(39) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state7;
    assign seq_loop_intf_10.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.pre_loop_state1 = 39'h0;
    assign seq_loop_intf_10.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.pre_loop_state2 = 39'h0;
    assign seq_loop_intf_10.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state4;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 39'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.post_loop_state2 = 39'h0;
    assign seq_loop_intf_10.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_10.post_loop_state3 = 39'h0;
    assign seq_loop_intf_10.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state9;
    assign seq_loop_intf_10.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_10.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_10.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_10.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state8;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state13;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(39) seq_loop_monitor_10;
    seq_loop_intf#(39) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state3;
    assign seq_loop_intf_11.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.pre_loop_state1 = 39'h0;
    assign seq_loop_intf_11.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.pre_loop_state2 = 39'h0;
    assign seq_loop_intf_11.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state14;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state17;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_11.post_loop_state2 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state34;
    assign seq_loop_intf_11.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_11.post_loop_state3 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state35;
    assign seq_loop_intf_11.post_states_valid[3] = 1'b1;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state4;
    assign seq_loop_intf_11.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_11.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_11.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_11.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state4;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state9;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(39) seq_loop_monitor_11;
    seq_loop_intf#(39) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state35;
    assign seq_loop_intf_12.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.pre_loop_state1 = 39'h0;
    assign seq_loop_intf_12.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.pre_loop_state2 = 39'h0;
    assign seq_loop_intf_12.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state25;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = 39'h0;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.post_loop_state2 = 39'h0;
    assign seq_loop_intf_12.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_12.post_loop_state3 = 39'h0;
    assign seq_loop_intf_12.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state36;
    assign seq_loop_intf_12.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_12.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_12.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_12.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state36;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state39;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(39) seq_loop_monitor_12;
    seq_loop_intf#(39) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state30;
    assign seq_loop_intf_13.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.pre_loop_state1 = 39'h0;
    assign seq_loop_intf_13.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.pre_loop_state2 = 39'h0;
    assign seq_loop_intf_13.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state25;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = 39'h0;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.post_loop_state2 = 39'h0;
    assign seq_loop_intf_13.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_13.post_loop_state3 = 39'h0;
    assign seq_loop_intf_13.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state31;
    assign seq_loop_intf_13.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_13.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_13.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_13.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state31;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state33;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(39) seq_loop_monitor_13;
    seq_loop_intf#(39) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state20;
    assign seq_loop_intf_14.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.pre_loop_state1 = 39'h0;
    assign seq_loop_intf_14.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.pre_loop_state2 = 39'h0;
    assign seq_loop_intf_14.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state25;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = 39'h0;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.post_loop_state2 = 39'h0;
    assign seq_loop_intf_14.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_14.post_loop_state3 = 39'h0;
    assign seq_loop_intf_14.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state24;
    assign seq_loop_intf_14.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_14.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_14.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_14.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state21;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state24;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(39) seq_loop_monitor_14;
    seq_loop_intf#(39) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state24;
    assign seq_loop_intf_15.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.pre_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state31;
    assign seq_loop_intf_15.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_15.pre_loop_state2 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state36;
    assign seq_loop_intf_15.pre_states_valid[2] = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state1;
    assign seq_loop_intf_15.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.post_loop_state1 = 39'h0;
    assign seq_loop_intf_15.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.post_loop_state2 = 39'h0;
    assign seq_loop_intf_15.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_15.post_loop_state3 = 39'h0;
    assign seq_loop_intf_15.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state25;
    assign seq_loop_intf_15.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.quit_loop_state1 = 39'h0;
    assign seq_loop_intf_15.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state2 = 39'h0;
    assign seq_loop_intf_15.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_15.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state25;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.ap_ST_fsm_state28;
    assign seq_loop_intf_15.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(39) seq_loop_monitor_15;
    seq_loop_intf#(5) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state1;
    assign seq_loop_intf_16.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_16.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_16.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state4;
    assign seq_loop_intf_16.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state5;
    assign seq_loop_intf_16.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_16.post_loop_state2 = 5'h0;
    assign seq_loop_intf_16.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_16.post_loop_state3 = 5'h0;
    assign seq_loop_intf_16.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state3;
    assign seq_loop_intf_16.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_16.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_16.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_16.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state2;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_377_1_fu_473.ap_ST_fsm_state3;
    assign seq_loop_intf_16.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(5) seq_loop_monitor_16;
    seq_loop_intf#(57) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state15;
    assign seq_loop_intf_17.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.pre_loop_state1 = 57'h0;
    assign seq_loop_intf_17.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.pre_loop_state2 = 57'h0;
    assign seq_loop_intf_17.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state52;
    assign seq_loop_intf_17.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state41;
    assign seq_loop_intf_17.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_17.post_loop_state2 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state23;
    assign seq_loop_intf_17.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_17.post_loop_state3 = 57'h0;
    assign seq_loop_intf_17.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state16;
    assign seq_loop_intf_17.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.quit_loop_state1 = 57'h0;
    assign seq_loop_intf_17.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state2 = 57'h0;
    assign seq_loop_intf_17.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_17.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state16;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state22;
    assign seq_loop_intf_17.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_17.one_state_loop = 1'b0;
    assign seq_loop_intf_17.one_state_block = 1'b0;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(57) seq_loop_monitor_17;
    seq_loop_intf#(57) seq_loop_intf_18(clock,reset);
    assign seq_loop_intf_18.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state31;
    assign seq_loop_intf_18.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.pre_loop_state1 = 57'h0;
    assign seq_loop_intf_18.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.pre_loop_state2 = 57'h0;
    assign seq_loop_intf_18.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_18.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state57;
    assign seq_loop_intf_18.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state23;
    assign seq_loop_intf_18.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_18.post_loop_state2 = 57'h0;
    assign seq_loop_intf_18.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_18.post_loop_state3 = 57'h0;
    assign seq_loop_intf_18.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_18.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state33;
    assign seq_loop_intf_18.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.quit_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state40;
    assign seq_loop_intf_18.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_18.quit_loop_state2 = 57'h0;
    assign seq_loop_intf_18.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_18.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_CS_fsm;
    assign seq_loop_intf_18.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state32;
    assign seq_loop_intf_18.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state40;
    assign seq_loop_intf_18.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_18.one_state_loop = 1'b0;
    assign seq_loop_intf_18.one_state_block = 1'b0;
    assign seq_loop_intf_18.finish = finish;
    csv_file_dump seq_loop_csv_dumper_18;
    seq_loop_monitor #(57) seq_loop_monitor_18;
    seq_loop_intf#(57) seq_loop_intf_19(clock,reset);
    assign seq_loop_intf_19.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state16;
    assign seq_loop_intf_19.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.pre_loop_state1 = 57'h0;
    assign seq_loop_intf_19.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.pre_loop_state2 = 57'h0;
    assign seq_loop_intf_19.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_19.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state41;
    assign seq_loop_intf_19.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state57;
    assign seq_loop_intf_19.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_19.post_loop_state2 = 57'h0;
    assign seq_loop_intf_19.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_19.post_loop_state3 = 57'h0;
    assign seq_loop_intf_19.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_19.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state23;
    assign seq_loop_intf_19.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.quit_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state33;
    assign seq_loop_intf_19.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_19.quit_loop_state2 = 57'h0;
    assign seq_loop_intf_19.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_19.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_CS_fsm;
    assign seq_loop_intf_19.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state23;
    assign seq_loop_intf_19.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state40;
    assign seq_loop_intf_19.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_19.one_state_loop = 1'b0;
    assign seq_loop_intf_19.one_state_block = 1'b0;
    assign seq_loop_intf_19.finish = finish;
    csv_file_dump seq_loop_csv_dumper_19;
    seq_loop_monitor #(57) seq_loop_monitor_19;
    seq_loop_intf#(57) seq_loop_intf_20(clock,reset);
    assign seq_loop_intf_20.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state12;
    assign seq_loop_intf_20.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.pre_loop_state1 = 57'h0;
    assign seq_loop_intf_20.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.pre_loop_state2 = 57'h0;
    assign seq_loop_intf_20.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_20.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state57;
    assign seq_loop_intf_20.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.post_loop_state1 = 57'h0;
    assign seq_loop_intf_20.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.post_loop_state2 = 57'h0;
    assign seq_loop_intf_20.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_20.post_loop_state3 = 57'h0;
    assign seq_loop_intf_20.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_20.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state13;
    assign seq_loop_intf_20.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.quit_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state33;
    assign seq_loop_intf_20.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_20.quit_loop_state2 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state55;
    assign seq_loop_intf_20.quit_states_valid[2] = 1'b1;
    assign seq_loop_intf_20.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_CS_fsm;
    assign seq_loop_intf_20.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state13;
    assign seq_loop_intf_20.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.ap_ST_fsm_state55;
    assign seq_loop_intf_20.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_20.one_state_loop = 1'b0;
    assign seq_loop_intf_20.one_state_block = 1'b0;
    assign seq_loop_intf_20.finish = finish;
    csv_file_dump seq_loop_csv_dumper_20;
    seq_loop_monitor #(57) seq_loop_monitor_20;
    seq_loop_intf#(5) seq_loop_intf_21(clock,reset);
    assign seq_loop_intf_21.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state1;
    assign seq_loop_intf_21.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_21.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_21.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_21.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state4;
    assign seq_loop_intf_21.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state5;
    assign seq_loop_intf_21.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_21.post_loop_state2 = 5'h0;
    assign seq_loop_intf_21.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_21.post_loop_state3 = 5'h0;
    assign seq_loop_intf_21.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_21.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state3;
    assign seq_loop_intf_21.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_21.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_21.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_21.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_CS_fsm;
    assign seq_loop_intf_21.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state2;
    assign seq_loop_intf_21.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_14_1_fu_587.ap_ST_fsm_state3;
    assign seq_loop_intf_21.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_21.one_state_loop = 1'b0;
    assign seq_loop_intf_21.one_state_block = 1'b0;
    assign seq_loop_intf_21.finish = finish;
    csv_file_dump seq_loop_csv_dumper_21;
    seq_loop_monitor #(5) seq_loop_monitor_21;
    seq_loop_intf#(5) seq_loop_intf_22(clock,reset);
    assign seq_loop_intf_22.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state1;
    assign seq_loop_intf_22.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_22.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_22.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_22.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state4;
    assign seq_loop_intf_22.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state5;
    assign seq_loop_intf_22.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_22.post_loop_state2 = 5'h0;
    assign seq_loop_intf_22.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_22.post_loop_state3 = 5'h0;
    assign seq_loop_intf_22.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_22.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state3;
    assign seq_loop_intf_22.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_22.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_22.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_22.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_CS_fsm;
    assign seq_loop_intf_22.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state2;
    assign seq_loop_intf_22.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_32_1_fu_596.ap_ST_fsm_state3;
    assign seq_loop_intf_22.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_22.one_state_loop = 1'b0;
    assign seq_loop_intf_22.one_state_block = 1'b0;
    assign seq_loop_intf_22.finish = finish;
    csv_file_dump seq_loop_csv_dumper_22;
    seq_loop_monitor #(5) seq_loop_monitor_22;
    seq_loop_intf#(5) seq_loop_intf_23(clock,reset);
    assign seq_loop_intf_23.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state1;
    assign seq_loop_intf_23.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_23.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_23.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_23.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state4;
    assign seq_loop_intf_23.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state5;
    assign seq_loop_intf_23.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_23.post_loop_state2 = 5'h0;
    assign seq_loop_intf_23.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_23.post_loop_state3 = 5'h0;
    assign seq_loop_intf_23.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_23.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state3;
    assign seq_loop_intf_23.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_23.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_23.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_23.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_CS_fsm;
    assign seq_loop_intf_23.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state2;
    assign seq_loop_intf_23.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_39_2_fu_606.ap_ST_fsm_state3;
    assign seq_loop_intf_23.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_23.one_state_loop = 1'b0;
    assign seq_loop_intf_23.one_state_block = 1'b0;
    assign seq_loop_intf_23.finish = finish;
    csv_file_dump seq_loop_csv_dumper_23;
    seq_loop_monitor #(5) seq_loop_monitor_23;
    seq_loop_intf#(5) seq_loop_intf_24(clock,reset);
    assign seq_loop_intf_24.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state1;
    assign seq_loop_intf_24.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_24.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_24.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_24.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state4;
    assign seq_loop_intf_24.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state5;
    assign seq_loop_intf_24.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_24.post_loop_state2 = 5'h0;
    assign seq_loop_intf_24.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_24.post_loop_state3 = 5'h0;
    assign seq_loop_intf_24.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_24.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state3;
    assign seq_loop_intf_24.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_24.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_24.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_24.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_CS_fsm;
    assign seq_loop_intf_24.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state2;
    assign seq_loop_intf_24.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_188_1_fu_365.ap_ST_fsm_state3;
    assign seq_loop_intf_24.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_24.one_state_loop = 1'b0;
    assign seq_loop_intf_24.one_state_block = 1'b0;
    assign seq_loop_intf_24.finish = finish;
    csv_file_dump seq_loop_csv_dumper_24;
    seq_loop_monitor #(5) seq_loop_monitor_24;
    seq_loop_intf#(7) seq_loop_intf_25(clock,reset);
    assign seq_loop_intf_25.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state1;
    assign seq_loop_intf_25.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_25.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.pre_loop_state2 = 7'h0;
    assign seq_loop_intf_25.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_25.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state6;
    assign seq_loop_intf_25.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state7;
    assign seq_loop_intf_25.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_25.post_loop_state2 = 7'h0;
    assign seq_loop_intf_25.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_25.post_loop_state3 = 7'h0;
    assign seq_loop_intf_25.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_25.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state5;
    assign seq_loop_intf_25.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_25.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.quit_loop_state2 = 7'h0;
    assign seq_loop_intf_25.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_25.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_CS_fsm;
    assign seq_loop_intf_25.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state2;
    assign seq_loop_intf_25.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_199_2_VITIS_LOOP_233_3_fu_373.ap_ST_fsm_state5;
    assign seq_loop_intf_25.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_25.one_state_loop = 1'b0;
    assign seq_loop_intf_25.one_state_block = 1'b0;
    assign seq_loop_intf_25.finish = finish;
    csv_file_dump seq_loop_csv_dumper_25;
    seq_loop_monitor #(7) seq_loop_monitor_25;
    seq_loop_intf#(5) seq_loop_intf_26(clock,reset);
    assign seq_loop_intf_26.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state1;
    assign seq_loop_intf_26.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_26.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_26.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_26.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state4;
    assign seq_loop_intf_26.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state5;
    assign seq_loop_intf_26.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_26.post_loop_state2 = 5'h0;
    assign seq_loop_intf_26.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_26.post_loop_state3 = 5'h0;
    assign seq_loop_intf_26.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_26.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state3;
    assign seq_loop_intf_26.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_26.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_26.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_26.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_CS_fsm;
    assign seq_loop_intf_26.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state2;
    assign seq_loop_intf_26.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_53_1_fu_168.ap_ST_fsm_state3;
    assign seq_loop_intf_26.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_26.one_state_loop = 1'b0;
    assign seq_loop_intf_26.one_state_block = 1'b0;
    assign seq_loop_intf_26.finish = finish;
    csv_file_dump seq_loop_csv_dumper_26;
    seq_loop_monitor #(5) seq_loop_monitor_26;
    seq_loop_intf#(5) seq_loop_intf_27(clock,reset);
    assign seq_loop_intf_27.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state1;
    assign seq_loop_intf_27.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_27.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_27.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_27.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state4;
    assign seq_loop_intf_27.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state5;
    assign seq_loop_intf_27.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_27.post_loop_state2 = 5'h0;
    assign seq_loop_intf_27.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_27.post_loop_state3 = 5'h0;
    assign seq_loop_intf_27.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_27.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state3;
    assign seq_loop_intf_27.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_27.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_27.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_27.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_CS_fsm;
    assign seq_loop_intf_27.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state2;
    assign seq_loop_intf_27.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_61_2_fu_176.ap_ST_fsm_state3;
    assign seq_loop_intf_27.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_27.one_state_loop = 1'b0;
    assign seq_loop_intf_27.one_state_block = 1'b0;
    assign seq_loop_intf_27.finish = finish;
    csv_file_dump seq_loop_csv_dumper_27;
    seq_loop_monitor #(5) seq_loop_monitor_27;
    seq_loop_intf#(5) seq_loop_intf_28(clock,reset);
    assign seq_loop_intf_28.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state1;
    assign seq_loop_intf_28.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_28.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_28.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_28.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state4;
    assign seq_loop_intf_28.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state5;
    assign seq_loop_intf_28.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_28.post_loop_state2 = 5'h0;
    assign seq_loop_intf_28.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_28.post_loop_state3 = 5'h0;
    assign seq_loop_intf_28.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_28.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state3;
    assign seq_loop_intf_28.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_28.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_28.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_28.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_CS_fsm;
    assign seq_loop_intf_28.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state2;
    assign seq_loop_intf_28.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_69_3_fu_185.ap_ST_fsm_state3;
    assign seq_loop_intf_28.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_28.one_state_loop = 1'b0;
    assign seq_loop_intf_28.one_state_block = 1'b0;
    assign seq_loop_intf_28.finish = finish;
    csv_file_dump seq_loop_csv_dumper_28;
    seq_loop_monitor #(5) seq_loop_monitor_28;
    seq_loop_intf#(5) seq_loop_intf_29(clock,reset);
    assign seq_loop_intf_29.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state1;
    assign seq_loop_intf_29.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_29.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_29.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_29.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state4;
    assign seq_loop_intf_29.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state5;
    assign seq_loop_intf_29.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_29.post_loop_state2 = 5'h0;
    assign seq_loop_intf_29.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_29.post_loop_state3 = 5'h0;
    assign seq_loop_intf_29.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_29.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state3;
    assign seq_loop_intf_29.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_29.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_29.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_29.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_CS_fsm;
    assign seq_loop_intf_29.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state2;
    assign seq_loop_intf_29.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_75_4_fu_193.ap_ST_fsm_state3;
    assign seq_loop_intf_29.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_29.one_state_loop = 1'b0;
    assign seq_loop_intf_29.one_state_block = 1'b0;
    assign seq_loop_intf_29.finish = finish;
    csv_file_dump seq_loop_csv_dumper_29;
    seq_loop_monitor #(5) seq_loop_monitor_29;
    seq_loop_intf#(5) seq_loop_intf_30(clock,reset);
    assign seq_loop_intf_30.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state1;
    assign seq_loop_intf_30.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_30.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_30.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_30.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state4;
    assign seq_loop_intf_30.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state5;
    assign seq_loop_intf_30.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_30.post_loop_state2 = 5'h0;
    assign seq_loop_intf_30.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_30.post_loop_state3 = 5'h0;
    assign seq_loop_intf_30.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_30.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state3;
    assign seq_loop_intf_30.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_30.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_30.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_30.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_CS_fsm;
    assign seq_loop_intf_30.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state2;
    assign seq_loop_intf_30.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_83_5_fu_201.ap_ST_fsm_state3;
    assign seq_loop_intf_30.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_30.one_state_loop = 1'b0;
    assign seq_loop_intf_30.one_state_block = 1'b0;
    assign seq_loop_intf_30.finish = finish;
    csv_file_dump seq_loop_csv_dumper_30;
    seq_loop_monitor #(5) seq_loop_monitor_30;
    seq_loop_intf#(5) seq_loop_intf_31(clock,reset);
    assign seq_loop_intf_31.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state1;
    assign seq_loop_intf_31.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_31.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_31.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_31.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state4;
    assign seq_loop_intf_31.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state5;
    assign seq_loop_intf_31.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_31.post_loop_state2 = 5'h0;
    assign seq_loop_intf_31.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_31.post_loop_state3 = 5'h0;
    assign seq_loop_intf_31.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_31.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state3;
    assign seq_loop_intf_31.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_31.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_31.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_31.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_CS_fsm;
    assign seq_loop_intf_31.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state2;
    assign seq_loop_intf_31.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_94_6_fu_210.ap_ST_fsm_state3;
    assign seq_loop_intf_31.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_31.one_state_loop = 1'b0;
    assign seq_loop_intf_31.one_state_block = 1'b0;
    assign seq_loop_intf_31.finish = finish;
    csv_file_dump seq_loop_csv_dumper_31;
    seq_loop_monitor #(5) seq_loop_monitor_31;
    seq_loop_intf#(5) seq_loop_intf_32(clock,reset);
    assign seq_loop_intf_32.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state1;
    assign seq_loop_intf_32.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_32.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_32.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_32.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state4;
    assign seq_loop_intf_32.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state5;
    assign seq_loop_intf_32.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_32.post_loop_state2 = 5'h0;
    assign seq_loop_intf_32.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_32.post_loop_state3 = 5'h0;
    assign seq_loop_intf_32.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_32.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state3;
    assign seq_loop_intf_32.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_32.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_32.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_32.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_CS_fsm;
    assign seq_loop_intf_32.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state2;
    assign seq_loop_intf_32.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_102_7_fu_219.ap_ST_fsm_state3;
    assign seq_loop_intf_32.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_32.one_state_loop = 1'b0;
    assign seq_loop_intf_32.one_state_block = 1'b0;
    assign seq_loop_intf_32.finish = finish;
    csv_file_dump seq_loop_csv_dumper_32;
    seq_loop_monitor #(5) seq_loop_monitor_32;
    seq_loop_intf#(5) seq_loop_intf_33(clock,reset);
    assign seq_loop_intf_33.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state1;
    assign seq_loop_intf_33.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_33.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_33.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_33.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state4;
    assign seq_loop_intf_33.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state5;
    assign seq_loop_intf_33.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_33.post_loop_state2 = 5'h0;
    assign seq_loop_intf_33.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_33.post_loop_state3 = 5'h0;
    assign seq_loop_intf_33.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_33.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state3;
    assign seq_loop_intf_33.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_33.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_33.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_33.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_CS_fsm;
    assign seq_loop_intf_33.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state2;
    assign seq_loop_intf_33.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_108_8_fu_227.ap_ST_fsm_state3;
    assign seq_loop_intf_33.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_33.one_state_loop = 1'b0;
    assign seq_loop_intf_33.one_state_block = 1'b0;
    assign seq_loop_intf_33.finish = finish;
    csv_file_dump seq_loop_csv_dumper_33;
    seq_loop_monitor #(5) seq_loop_monitor_33;
    seq_loop_intf#(5) seq_loop_intf_34(clock,reset);
    assign seq_loop_intf_34.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state1;
    assign seq_loop_intf_34.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_34.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_34.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_34.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state4;
    assign seq_loop_intf_34.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state5;
    assign seq_loop_intf_34.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_34.post_loop_state2 = 5'h0;
    assign seq_loop_intf_34.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_34.post_loop_state3 = 5'h0;
    assign seq_loop_intf_34.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_34.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state3;
    assign seq_loop_intf_34.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_34.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_34.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_34.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_CS_fsm;
    assign seq_loop_intf_34.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state2;
    assign seq_loop_intf_34.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_Dependency_Update_BypassMode_SrcTgt_fu_667.grp_Dependency_Update_BypassMode_SrcTgt_Pipeline_VITIS_LOOP_116_9_fu_235.ap_ST_fsm_state3;
    assign seq_loop_intf_34.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_34.one_state_loop = 1'b0;
    assign seq_loop_intf_34.one_state_block = 1'b0;
    assign seq_loop_intf_34.finish = finish;
    csv_file_dump seq_loop_csv_dumper_34;
    seq_loop_monitor #(5) seq_loop_monitor_34;
    seq_loop_intf#(5) seq_loop_intf_35(clock,reset);
    assign seq_loop_intf_35.pre_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state1;
    assign seq_loop_intf_35.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.pre_loop_state1 = 5'h0;
    assign seq_loop_intf_35.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.pre_loop_state2 = 5'h0;
    assign seq_loop_intf_35.pre_states_valid[2] = 1'b0;
    assign seq_loop_intf_35.post_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state4;
    assign seq_loop_intf_35.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.post_loop_state1 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state5;
    assign seq_loop_intf_35.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_35.post_loop_state2 = 5'h0;
    assign seq_loop_intf_35.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_35.post_loop_state3 = 5'h0;
    assign seq_loop_intf_35.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_35.quit_loop_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state3;
    assign seq_loop_intf_35.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.quit_loop_state1 = 5'h0;
    assign seq_loop_intf_35.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.quit_loop_state2 = 5'h0;
    assign seq_loop_intf_35.quit_states_valid[2] = 1'b0;
    assign seq_loop_intf_35.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_CS_fsm;
    assign seq_loop_intf_35.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state2;
    assign seq_loop_intf_35.iter_end_state0 = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_RoutingAvailability_CheckPredecessor_and_Placement_Pipeline_VITIS_LOOP_127_1_fu_691.ap_ST_fsm_state3;
    assign seq_loop_intf_35.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_35.one_state_loop = 1'b0;
    assign seq_loop_intf_35.one_state_block = 1'b0;
    assign seq_loop_intf_35.finish = finish;
    csv_file_dump seq_loop_csv_dumper_35;
    seq_loop_monitor #(5) seq_loop_monitor_35;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_1.quit_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_1.loop_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_685_5_VITIS_LOOP_686_6_VITIS_LOOP_687_7_fu_191.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.quit_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.loop_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_697_10_VITIS_LOOP_698_11_VITIS_LOOP_699_12_fu_203.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b0;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_3.quit_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_3.loop_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_724_19_VITIS_LOOP_726_20_fu_239.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_4.quit_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_enable_reg_pp0_iter3;
    assign upc_loop_intf_4.loop_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_736_21_VITIS_LOOP_738_22_fu_249.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.loop_start = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_runOne.grp_Reset_fu_334.grp_Reset_Pipeline_VITIS_LOOP_719_18_fu_259.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b0;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_470_5_fu_522.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_497_8_VITIS_LOOP_498_9_fu_540.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b0;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_508_10_fu_551.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b0;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_CurOptPotentialPlacement_List_BypassLess_Gen_fu_439.grp_CurOptPotentialPlacement_List_BypassLess_Gen_Pipeline_VITIS_LOOP_562_14_fu_559.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b0;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_398_3_fu_493.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b0;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(2) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_RoutingAvailability_CheckPredecessor_and_Placement_fu_507.grp_BypassOptPlacement_Gen_Record_fu_615.grp_BypassOptPlacement_Gen_Record_Pipeline_VITIS_LOOP_255_5_fu_420.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(2) upc_loop_monitor_11;
    upc_loop_intf#(1) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.loop_start = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_runOne.grp_dynamic_placement_routing_fu_400.grp_dynamic_placement_routing_Pipeline_VITIS_LOOP_415_5_fu_597.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b0;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(1) upc_loop_monitor_12;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);
    seq_loop_csv_dumper_18 = new("./seq_loop_status18.csv");
    seq_loop_monitor_18 = new(seq_loop_intf_18,seq_loop_csv_dumper_18);
    seq_loop_csv_dumper_19 = new("./seq_loop_status19.csv");
    seq_loop_monitor_19 = new(seq_loop_intf_19,seq_loop_csv_dumper_19);
    seq_loop_csv_dumper_20 = new("./seq_loop_status20.csv");
    seq_loop_monitor_20 = new(seq_loop_intf_20,seq_loop_csv_dumper_20);
    seq_loop_csv_dumper_21 = new("./seq_loop_status21.csv");
    seq_loop_monitor_21 = new(seq_loop_intf_21,seq_loop_csv_dumper_21);
    seq_loop_csv_dumper_22 = new("./seq_loop_status22.csv");
    seq_loop_monitor_22 = new(seq_loop_intf_22,seq_loop_csv_dumper_22);
    seq_loop_csv_dumper_23 = new("./seq_loop_status23.csv");
    seq_loop_monitor_23 = new(seq_loop_intf_23,seq_loop_csv_dumper_23);
    seq_loop_csv_dumper_24 = new("./seq_loop_status24.csv");
    seq_loop_monitor_24 = new(seq_loop_intf_24,seq_loop_csv_dumper_24);
    seq_loop_csv_dumper_25 = new("./seq_loop_status25.csv");
    seq_loop_monitor_25 = new(seq_loop_intf_25,seq_loop_csv_dumper_25);
    seq_loop_csv_dumper_26 = new("./seq_loop_status26.csv");
    seq_loop_monitor_26 = new(seq_loop_intf_26,seq_loop_csv_dumper_26);
    seq_loop_csv_dumper_27 = new("./seq_loop_status27.csv");
    seq_loop_monitor_27 = new(seq_loop_intf_27,seq_loop_csv_dumper_27);
    seq_loop_csv_dumper_28 = new("./seq_loop_status28.csv");
    seq_loop_monitor_28 = new(seq_loop_intf_28,seq_loop_csv_dumper_28);
    seq_loop_csv_dumper_29 = new("./seq_loop_status29.csv");
    seq_loop_monitor_29 = new(seq_loop_intf_29,seq_loop_csv_dumper_29);
    seq_loop_csv_dumper_30 = new("./seq_loop_status30.csv");
    seq_loop_monitor_30 = new(seq_loop_intf_30,seq_loop_csv_dumper_30);
    seq_loop_csv_dumper_31 = new("./seq_loop_status31.csv");
    seq_loop_monitor_31 = new(seq_loop_intf_31,seq_loop_csv_dumper_31);
    seq_loop_csv_dumper_32 = new("./seq_loop_status32.csv");
    seq_loop_monitor_32 = new(seq_loop_intf_32,seq_loop_csv_dumper_32);
    seq_loop_csv_dumper_33 = new("./seq_loop_status33.csv");
    seq_loop_monitor_33 = new(seq_loop_intf_33,seq_loop_csv_dumper_33);
    seq_loop_csv_dumper_34 = new("./seq_loop_status34.csv");
    seq_loop_monitor_34 = new(seq_loop_intf_34,seq_loop_csv_dumper_34);
    seq_loop_csv_dumper_35 = new("./seq_loop_status35.csv");
    seq_loop_monitor_35 = new(seq_loop_intf_35,seq_loop_csv_dumper_35);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_19);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_20);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_21);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_22);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_23);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_24);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_25);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_26);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_27);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_28);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_29);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_30);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_31);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_32);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_33);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_34);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_35);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
